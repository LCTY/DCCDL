module main(
    );

	
	dff s0(Clk, Reset, LdEnable, d_0, Load, q_0);
	dff s1(Clk, Reset, LdEnable, d_1, Load, q_1);
	dff s2(Clk, Reset, LdEnable, q_0, Load, q_2);
	
	xor ()
	
	xor 

endmodule
